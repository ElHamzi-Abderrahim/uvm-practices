`ifndef MD_PKG_SV
`define MD_PKG_SV

    `include "md_if.sv"

    package md_pkg ;
        import uvm_pkg::* ;

        `include "md_reset_handler.sv"
        
        `include "md_item_base.sv"
        `include "md_item_drv.sv"
        `include "md_item_drv_master.sv"
        
        `include "md_agent_config.sv"
        `include "md_agent_config_slave.sv"
        `include "md_agent_config_master.sv"
        
        `include "md_sequencer.sv"
        `include "md_sequencer_master.sv"
        
        `include "md_driver.sv"
        `include "md_driver_master.sv"
        
        `include "md_agent.sv"
        `include "md_agent_slave.sv"
        `include "md_agent_master.sv"

        `include "md_sequence_base.sv"
        `include "md_sequence_simple_master.sv"


    endpackage

`endif