`ifndef TEST_DEFINES_SV
`define TEST_DEFINES_SV

    `ifndef ALIGN_TEST_DATA_WIDTH
        `define ALIGN_TEST_DATA_WIDTH 32
    `endif


`endif
