`ifndef APB_TYPES_SV
  	`define APB_TYPES_SV
	
	// Virtual interface type:
	typedef virtual apb_if apb_vif;
	
`endif